module code;
    initial begin $display("Hello World"); $finish; end
endmodule
